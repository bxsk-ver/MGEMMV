module GP_Gen_1_49 #(
    parameter width=49
)( 
    input wire [width:1] p,
    input wire [width:1] g,
    output wire [width:1] P,
    output wire [width:1] G
);
    wire p_33_49, p_33_48, p_33_47, p_33_46, p_33_45, p_33_44, p_33_43, p_33_42, p_33_41, p_33_40, p_33_39, p_33_38, p_33_37, p_33_36, p_33_35, p_33_34, p_33_33;
    wire g_33_49, g_33_48, g_33_47, g_33_46, g_33_45, g_33_44, g_33_43, g_33_42, g_33_41, g_33_40, g_33_39, g_33_38, g_33_37, g_33_36, g_33_35, g_33_34, g_33_33;
    GP_Gen_1_32 #(.width(32)) u0 (.p(p[32:1]), .g(g[32:1]), .P(P[32:1]), .G(G[32:1]));
    GP_Gen_1_17 #(.width(17)) u1 (.p(p[49:33]), .g(g[49:33]), .P({p_33_49, p_33_48, p_33_47, p_33_46, p_33_45, p_33_44, p_33_43, p_33_42, p_33_41, p_33_40, p_33_39, p_33_38, p_33_37, p_33_36, p_33_35, p_33_34, p_33_33}), .G({g_33_49, g_33_48, g_33_47, g_33_46, g_33_45, g_33_44, g_33_43, g_33_42, g_33_41, g_33_40, g_33_39, g_33_38, g_33_37, g_33_36, g_33_35, g_33_34, g_33_33}));
    assign P[33] = P[32] & p_33_33;
    assign G[33] = g_33_33 | (G[32] & p_33_33);
    assign P[34] = P[32] & p_33_34;
    assign G[34] = g_33_34 | (G[32] & p_33_34);
    assign P[35] = P[32] & p_33_35;
    assign G[35] = g_33_35 | (G[32] & p_33_35);
    assign P[36] = P[32] & p_33_36;
    assign G[36] = g_33_36 | (G[32] & p_33_36);
    assign P[37] = P[32] & p_33_37;
    assign G[37] = g_33_37 | (G[32] & p_33_37);
    assign P[38] = P[32] & p_33_38;
    assign G[38] = g_33_38 | (G[32] & p_33_38);
    assign P[39] = P[32] & p_33_39;
    assign G[39] = g_33_39 | (G[32] & p_33_39);
    assign P[40] = P[32] & p_33_40;
    assign G[40] = g_33_40 | (G[32] & p_33_40);
    assign P[41] = P[32] & p_33_41;
    assign G[41] = g_33_41 | (G[32] & p_33_41);
    assign P[42] = P[32] & p_33_42;
    assign G[42] = g_33_42 | (G[32] & p_33_42);
    assign P[43] = P[32] & p_33_43;
    assign G[43] = g_33_43 | (G[32] & p_33_43);
    assign P[44] = P[32] & p_33_44;
    assign G[44] = g_33_44 | (G[32] & p_33_44);
    assign P[45] = P[32] & p_33_45;
    assign G[45] = g_33_45 | (G[32] & p_33_45);
    assign P[46] = P[32] & p_33_46;
    assign G[46] = g_33_46 | (G[32] & p_33_46);
    assign P[47] = P[32] & p_33_47;
    assign G[47] = g_33_47 | (G[32] & p_33_47);
    assign P[48] = P[32] & p_33_48;
    assign G[48] = g_33_48 | (G[32] & p_33_48);
    assign P[49] = P[32] & p_33_49;
    assign G[49] = g_33_49 | (G[32] & p_33_49);

endmodule
